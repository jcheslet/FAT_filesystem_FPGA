----------------------------------------------------------------------------------------------------
-- SDcard_raw_access_v2
----------------------------------------------------------------------------------------------------
