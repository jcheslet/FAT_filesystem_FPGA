----------------------------------------------------------------------------------
-- 
----------------------------------------------------------------------------------
