----------------------------------------------------------------------------------
-- Sdcard_readstream
----------------------------------------------------------------------------------
