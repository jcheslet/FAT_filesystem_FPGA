----------------------------------------------------------------------------------
-- SDcard_raw_access_simmodel
----------------------------------------------------------------------------------
