----------------------------------------------------------------------------------
-- Sdcard_writestream
----------------------------------------------------------------------------------
